
***** Spice Netlist for Cell 'Lab11_inv' *****

************** Module Lab11_inv **************
.subckt Lab11_inv NULL vin vout
m2 vout vin vdd vdd scmosp w='0.6u' l='0.4u' m='1' 
m1 vout vin gnd gnd scmosn w='0.6u' l='0.4u' m='1' 
.ends Lab11_inv




